library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VGA_sampler is
	port(
		clk_200M_i 		: in  std_logic	
	);
end VGA_sampler;

architecture Behavioral of VGA_sampler is

begin


end Behavioral;

