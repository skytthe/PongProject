library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package components is
		
end package components;

package body components is
	
end package body components;
