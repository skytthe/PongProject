library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity filter is
	port(
		clk_200M_i 		: in  std_logic	
	);
end filter;

architecture Behavioral of filter is

begin


end Behavioral;

