library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity graphics_engine is
	port(
		clk_200M_i 		: in  std_logic	
	);
end graphics_engine;

architecture Behavioral of graphics_engine is

begin


end Behavioral;

