library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity delay_chain is
end delay_chain;

architecture Behavioral of delay_chain is

begin


end Behavioral;

